`timescale 1ns/10ps

//   misc.v
//
//   Copyright 2024 Brady Etz
//
//   Licensed under the Apache License, Version 2.0 (the "License");
//   you may not use this file except in compliance with the License.
//   You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in writing, software
//   distributed under the License is distributed on an "AS IS" BASIS,
//   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//   See the License for the specific language governing permissions and
//   limitations under the License.


module clkdiv_by_2 (
  input      clk_i, rstn_i,
  output reg clk_o
);
  always @(posedge clk_i or negedge rstn_i) begin
    if (!rstn_i) clk_o <= 1'b0;
    else clk_o <= ~clk_o;
  end
endmodule


// Ripple counter stage with common clk_i
// Useful for FPGAs and tight setup constraints
module ripple_stage (
  input      clk_i, rstn_i,
  input      in,
  output reg out
);
  wire enable; reg in_r;
  assign enable = in & ~in_r;
  
  always @(posedge clk_i or negedge rstn_i) begin
    if (!rstn_i) begin
      in_r <= 1'b0; out <= 1'b0;
    end else begin
      in_r <= in;
      if (enable) out <= ~out;
    end
  end
endmodule
